`define numLayers 5
`define dataWidth 16
`define numNeuronLayer1 30
`define numWeightLayer1 784
`define Layer1ActType "relu"
`define numNeuronLayer2 30
`define numWeightLayer2 30
`define Layer2ActType "relu"
`define numNeuronLayer3 10
`define numWeightLayer3 30
`define Layer3ActType "relu"
`define numNeuronLayer4 10
`define numWeightLayer4 10
`define Layer4ActType "relu"
`define numNeuronLayer5 10
`define numWeightLayer5 10
`define Layer5ActType "hardmax"
`define sigmoidSize 5
`define weightIntWidth 4
`define WB_DIR "/home/huyld/WORK/neural_network/mnist/sim/training/w_b_correct/"
`define TEST_DIR "/home/huyld/WORK/neural_network/mnist/sim/training/testData/"
